interface intf();
  logic clk;
  logic rst;
  logic d;
  logic q;
endinterface
