interface inf;
  
  logic clk;
  logic rst;
  logic [3:0] count;
  
endinterface
